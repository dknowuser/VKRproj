module trapezoidal_filter (input clk);
endmodule